module out

pub fn print_some_thing() {
	println("You SUCKS, your d*ck")
}

pub fn i_dunno() {
	a := 50
	println("The value of a is {a}")
}