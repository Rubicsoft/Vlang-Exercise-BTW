module out

pub fn print_some_thing() {
	println("You SUCKS, your d*ck")
}